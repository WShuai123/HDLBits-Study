//使用一条 assign 语句，将输入端口的值赋给输出端口
module top_module( input in, output out );
	assign out=in;
endmodule
